module perceptron_top(
input logic                      clk,
input logic [ADDRESS_WIDTH-1:0]  pc,
input logic                      branch_result,



);



endmodule