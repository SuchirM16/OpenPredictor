module condition_checker
(

);


endmodule