
module weight_updater
(

);

endmodule